//This document contains test cases to verify snoop side behavior of L1 Cache
//Author : Abhishek Gupta

module multicore

//for verifying the fuctionality of muticore cache environment
