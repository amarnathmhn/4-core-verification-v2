import uvm_pkg::*;
`include "interfacesMultiCore.svh"
`include "uvm_macros.svh"
`include "helloworld.svh"
