	/*
	`include "cache_def_0.v"
	`include "cache_def_I_0.v"
	
	`include "cache_block_0.v" 
	`include "cache_block_1.v" 
	`include "cache_block_2.v" 
	`include "cache_block_3.v" 

	`include "cache_block_I_0.v" 
	`include "cache_block_I_1.v" 
	`include "cache_block_I_2.v" 
	`include "cache_block_I_3.v" 
	
	`include "cache_controller_0.v"
	`include "cache_controller_1.v"
	`include "cache_controller_2.v"
	`include "cache_controller_3.v"

	`include "cache_controller_I_0.v"
	`include "cache_controller_I_1.v"
	`include "cache_controller_I_2.v"
	`include "cache_controller_I_3.v"
	
	`include "cache_wrapper_0.v"
	`include "cache_wrapper_1.v"
	`include "cache_wrapper_2.v"
	`include "cache_wrapper_3.v"
	
	`include "cache_wrapper_I_0.v"
	`include "cache_wrapper_I_1.v"
	`include "cache_wrapper_I_2.v"
	`include "cache_wrapper_I_3.v"
*/
	
